`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:59:16 08/01/2018 
// Design Name: 
// Module Name:    ROMtest 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
//-- Fichero: genrom.v
module genrom #(           //-- Parametros
			parameter ROMFILE = "StageData.list",
         parameter AW = 9,   //-- Bits de las direcciones (Adress width)
         parameter DW = 32)   //-- Bits de los datos (Data witdh)

       (                              //-- Puertos
         input clk,                   //-- Se�al de reloj global
         input wire [AW-1: 0] addr,   //-- Direcciones
         output reg [DW-1: 0] data);  //-- Dato de salida

//-- Parametro: Nombre del fichero con el contenido de la ROM

//-- Calcular el numero de posiciones totales de memoria
localparam NPOS = 2 ** AW;

  //-- Memoria
  reg [DW-1: 0] rom [NPOS-1: 0];

  //-- Lectura de la memoria
  always @(posedge clk) begin
    data <= rom[addr];
  end

//-- Cargar en la memoria el fichero ROMFILE
//-- Los valores deben estan dados en hexadecimal
initial begin
  $readmemb(ROMFILE, rom);
end

endmodule
